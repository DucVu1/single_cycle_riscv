library verilog;
use verilog.vl_types.all;
entity barrel_shifter_right_32 is
    port(
        data            : in     vl_logic_vector(31 downto 0);
        type_shift      : in     vl_logic;
        amt             : in     vl_logic_vector(4 downto 0);
        \out\           : out    vl_logic_vector(31 downto 0)
    );
end barrel_shifter_right_32;
